module main

fn main() {
	println('Algorithms and data structures written in V language')
}
