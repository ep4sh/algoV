module main

fn main() {
	println('Algorythms and data structures written with V language')
}
