/*
* main.v
 * Copyright (C) 2021 Pasha Radchenko <ep4sh2k@gmail.com>
 *
 * Distributed under terms of the MIT license.
*/

module main

fn main() {
	println('Algorithms and data structures written in V language')
}
